//---------------------------------------------------------------------
// Title   : 1024x16 bit Sine wave dummy sample data
// Project : JESD204
//---------------------------------------------------------------------
// File    : sine16.vh
// Author  : Xilinx
//---------------------------------------------------------------------
// Description:
//
//---------------------------------------------------------------------
// (c) Copyright 2012-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
//
//----------------------------------------------------------------------------
  assign sine_lookup[0   ]    = 16'h8000;
  assign sine_lookup[1   ]    = 16'h80C9;
  assign sine_lookup[2   ]    = 16'h8192;
  assign sine_lookup[3   ]    = 16'h825B;
  assign sine_lookup[4   ]    = 16'h8324;
  assign sine_lookup[5   ]    = 16'h83ED;
  assign sine_lookup[6   ]    = 16'h84B6;
  assign sine_lookup[7   ]    = 16'h857F;
  assign sine_lookup[8   ]    = 16'h8648;
  assign sine_lookup[9   ]    = 16'h8711;
  assign sine_lookup[10  ]    = 16'h87D9;
  assign sine_lookup[11  ]    = 16'h88A2;
  assign sine_lookup[12  ]    = 16'h896A;
  assign sine_lookup[13  ]    = 16'h8A33;
  assign sine_lookup[14  ]    = 16'h8AFB;
  assign sine_lookup[15  ]    = 16'h8BC4;
  assign sine_lookup[16  ]    = 16'h8C8C;
  assign sine_lookup[17  ]    = 16'h8D54;
  assign sine_lookup[18  ]    = 16'h8E1C;
  assign sine_lookup[19  ]    = 16'h8EE3;
  assign sine_lookup[20  ]    = 16'h8FAB;
  assign sine_lookup[21  ]    = 16'h9072;
  assign sine_lookup[22  ]    = 16'h913A;
  assign sine_lookup[23  ]    = 16'h9201;
  assign sine_lookup[24  ]    = 16'h92C8;
  assign sine_lookup[25  ]    = 16'h938F;
  assign sine_lookup[26  ]    = 16'h9455;
  assign sine_lookup[27  ]    = 16'h951C;
  assign sine_lookup[28  ]    = 16'h95E2;
  assign sine_lookup[29  ]    = 16'h96A8;
  assign sine_lookup[30  ]    = 16'h976E;
  assign sine_lookup[31  ]    = 16'h9833;
  assign sine_lookup[32  ]    = 16'h98F9;
  assign sine_lookup[33  ]    = 16'h99BE;
  assign sine_lookup[34  ]    = 16'h9A82;
  assign sine_lookup[35  ]    = 16'h9B47;
  assign sine_lookup[36  ]    = 16'h9C0B;
  assign sine_lookup[37  ]    = 16'h9CCF;
  assign sine_lookup[38  ]    = 16'h9D93;
  assign sine_lookup[39  ]    = 16'h9E57;
  assign sine_lookup[40  ]    = 16'h9F1A;
  assign sine_lookup[41  ]    = 16'h9FDD;
  assign sine_lookup[42  ]    = 16'hA09F;
  assign sine_lookup[43  ]    = 16'hA161;
  assign sine_lookup[44  ]    = 16'hA223;
  assign sine_lookup[45  ]    = 16'hA2E5;
  assign sine_lookup[46  ]    = 16'hA3A6;
  assign sine_lookup[47  ]    = 16'hA467;
  assign sine_lookup[48  ]    = 16'hA528;
  assign sine_lookup[49  ]    = 16'hA5E8;
  assign sine_lookup[50  ]    = 16'hA6A8;
  assign sine_lookup[51  ]    = 16'hA767;
  assign sine_lookup[52  ]    = 16'hA826;
  assign sine_lookup[53  ]    = 16'hA8E5;
  assign sine_lookup[54  ]    = 16'hA9A3;
  assign sine_lookup[55  ]    = 16'hAA61;
  assign sine_lookup[56  ]    = 16'hAB1F;
  assign sine_lookup[57  ]    = 16'hABDC;
  assign sine_lookup[58  ]    = 16'hAC99;
  assign sine_lookup[59  ]    = 16'hAD55;
  assign sine_lookup[60  ]    = 16'hAE11;
  assign sine_lookup[61  ]    = 16'hAECC;
  assign sine_lookup[62  ]    = 16'hAF87;
  assign sine_lookup[63  ]    = 16'hB041;
  assign sine_lookup[64  ]    = 16'hB0FB;
  assign sine_lookup[65  ]    = 16'hB1B5;
  assign sine_lookup[66  ]    = 16'hB26E;
  assign sine_lookup[67  ]    = 16'hB326;
  assign sine_lookup[68  ]    = 16'hB3DF;
  assign sine_lookup[69  ]    = 16'hB496;
  assign sine_lookup[70  ]    = 16'hB54D;
  assign sine_lookup[71  ]    = 16'hB604;
  assign sine_lookup[72  ]    = 16'hB6BA;
  assign sine_lookup[73  ]    = 16'hB76F;
  assign sine_lookup[74  ]    = 16'hB824;
  assign sine_lookup[75  ]    = 16'hB8D9;
  assign sine_lookup[76  ]    = 16'hB98C;
  assign sine_lookup[77  ]    = 16'hBA40;
  assign sine_lookup[78  ]    = 16'hBAF2;
  assign sine_lookup[79  ]    = 16'hBBA5;
  assign sine_lookup[80  ]    = 16'hBC56;
  assign sine_lookup[81  ]    = 16'hBD07;
  assign sine_lookup[82  ]    = 16'hBDB8;
  assign sine_lookup[83  ]    = 16'hBE68;
  assign sine_lookup[84  ]    = 16'hBF17;
  assign sine_lookup[85  ]    = 16'hBFC5;
  assign sine_lookup[86  ]    = 16'hC073;
  assign sine_lookup[87  ]    = 16'hC121;
  assign sine_lookup[88  ]    = 16'hC1CE;
  assign sine_lookup[89  ]    = 16'hC27A;
  assign sine_lookup[90  ]    = 16'hC325;
  assign sine_lookup[91  ]    = 16'hC3D0;
  assign sine_lookup[92  ]    = 16'hC47A;
  assign sine_lookup[93  ]    = 16'hC524;
  assign sine_lookup[94  ]    = 16'hC5CD;
  assign sine_lookup[95  ]    = 16'hC675;
  assign sine_lookup[96  ]    = 16'hC71C;
  assign sine_lookup[97  ]    = 16'hC7C3;
  assign sine_lookup[98  ]    = 16'hC869;
  assign sine_lookup[99  ]    = 16'hC90F;
  assign sine_lookup[100 ]    = 16'hC9B4;
  assign sine_lookup[101 ]    = 16'hCA58;
  assign sine_lookup[102 ]    = 16'hCAFB;
  assign sine_lookup[103 ]    = 16'hCB9D;
  assign sine_lookup[104 ]    = 16'hCC3F;
  assign sine_lookup[105 ]    = 16'hCCE0;
  assign sine_lookup[106 ]    = 16'hCD81;
  assign sine_lookup[107 ]    = 16'hCE20;
  assign sine_lookup[108 ]    = 16'hCEBF;
  assign sine_lookup[109 ]    = 16'hCF5D;
  assign sine_lookup[110 ]    = 16'hCFFB;
  assign sine_lookup[111 ]    = 16'hD097;
  assign sine_lookup[112 ]    = 16'hD133;
  assign sine_lookup[113 ]    = 16'hD1CE;
  assign sine_lookup[114 ]    = 16'hD268;
  assign sine_lookup[115 ]    = 16'hD302;
  assign sine_lookup[116 ]    = 16'hD39B;
  assign sine_lookup[117 ]    = 16'hD432;
  assign sine_lookup[118 ]    = 16'hD4C9;
  assign sine_lookup[119 ]    = 16'hD560;
  assign sine_lookup[120 ]    = 16'hD5F5;
  assign sine_lookup[121 ]    = 16'hD68A;
  assign sine_lookup[122 ]    = 16'hD71D;
  assign sine_lookup[123 ]    = 16'hD7B0;
  assign sine_lookup[124 ]    = 16'hD842;
  assign sine_lookup[125 ]    = 16'hD8D3;
  assign sine_lookup[126 ]    = 16'hD964;
  assign sine_lookup[127 ]    = 16'hD9F3;
  assign sine_lookup[128 ]    = 16'hDA82;
  assign sine_lookup[129 ]    = 16'hDB0F;
  assign sine_lookup[130 ]    = 16'hDB9C;
  assign sine_lookup[131 ]    = 16'hDC28;
  assign sine_lookup[132 ]    = 16'hDCB3;
  assign sine_lookup[133 ]    = 16'hDD3E;
  assign sine_lookup[134 ]    = 16'hDDC7;
  assign sine_lookup[135 ]    = 16'hDE4F;
  assign sine_lookup[136 ]    = 16'hDED7;
  assign sine_lookup[137 ]    = 16'hDF5D;
  assign sine_lookup[138 ]    = 16'hDFE3;
  assign sine_lookup[139 ]    = 16'hE068;
  assign sine_lookup[140 ]    = 16'hE0EB;
  assign sine_lookup[141 ]    = 16'hE16E;
  assign sine_lookup[142 ]    = 16'hE1F0;
  assign sine_lookup[143 ]    = 16'hE271;
  assign sine_lookup[144 ]    = 16'hE2F1;
  assign sine_lookup[145 ]    = 16'hE370;
  assign sine_lookup[146 ]    = 16'hE3EE;
  assign sine_lookup[147 ]    = 16'hE46C;
  assign sine_lookup[148 ]    = 16'hE4E8;
  assign sine_lookup[149 ]    = 16'hE563;
  assign sine_lookup[150 ]    = 16'hE5DD;
  assign sine_lookup[151 ]    = 16'hE656;
  assign sine_lookup[152 ]    = 16'hE6CF;
  assign sine_lookup[153 ]    = 16'hE746;
  assign sine_lookup[154 ]    = 16'hE7BC;
  assign sine_lookup[155 ]    = 16'hE832;
  assign sine_lookup[156 ]    = 16'hE8A6;
  assign sine_lookup[157 ]    = 16'hE919;
  assign sine_lookup[158 ]    = 16'hE98B;
  assign sine_lookup[159 ]    = 16'hE9FD;
  assign sine_lookup[160 ]    = 16'hEA6D;
  assign sine_lookup[161 ]    = 16'hEADC;
  assign sine_lookup[162 ]    = 16'hEB4A;
  assign sine_lookup[163 ]    = 16'hEBB7;
  assign sine_lookup[164 ]    = 16'hEC23;
  assign sine_lookup[165 ]    = 16'hEC8E;
  assign sine_lookup[166 ]    = 16'hECF8;
  assign sine_lookup[167 ]    = 16'hED61;
  assign sine_lookup[168 ]    = 16'hEDC9;
  assign sine_lookup[169 ]    = 16'hEE30;
  assign sine_lookup[170 ]    = 16'hEE96;
  assign sine_lookup[171 ]    = 16'hEEFB;
  assign sine_lookup[172 ]    = 16'hEF5E;
  assign sine_lookup[173 ]    = 16'hEFC1;
  assign sine_lookup[174 ]    = 16'hF022;
  assign sine_lookup[175 ]    = 16'hF083;
  assign sine_lookup[176 ]    = 16'hF0E2;
  assign sine_lookup[177 ]    = 16'hF140;
  assign sine_lookup[178 ]    = 16'hF19D;
  assign sine_lookup[179 ]    = 16'hF1F9;
  assign sine_lookup[180 ]    = 16'hF254;
  assign sine_lookup[181 ]    = 16'hF2AE;
  assign sine_lookup[182 ]    = 16'hF307;
  assign sine_lookup[183 ]    = 16'hF35E;
  assign sine_lookup[184 ]    = 16'hF3B5;
  assign sine_lookup[185 ]    = 16'hF40A;
  assign sine_lookup[186 ]    = 16'hF45F;
  assign sine_lookup[187 ]    = 16'hF4B2;
  assign sine_lookup[188 ]    = 16'hF504;
  assign sine_lookup[189 ]    = 16'hF555;
  assign sine_lookup[190 ]    = 16'hF5A5;
  assign sine_lookup[191 ]    = 16'hF5F3;
  assign sine_lookup[192 ]    = 16'hF641;
  assign sine_lookup[193 ]    = 16'hF68D;
  assign sine_lookup[194 ]    = 16'hF6D8;
  assign sine_lookup[195 ]    = 16'hF722;
  assign sine_lookup[196 ]    = 16'hF76B;
  assign sine_lookup[197 ]    = 16'hF7B3;
  assign sine_lookup[198 ]    = 16'hF7FA;
  assign sine_lookup[199 ]    = 16'hF83F;
  assign sine_lookup[200 ]    = 16'hF884;
  assign sine_lookup[201 ]    = 16'hF8C7;
  assign sine_lookup[202 ]    = 16'hF909;
  assign sine_lookup[203 ]    = 16'hF94A;
  assign sine_lookup[204 ]    = 16'hF989;
  assign sine_lookup[205 ]    = 16'hF9C8;
  assign sine_lookup[206 ]    = 16'hFA05;
  assign sine_lookup[207 ]    = 16'hFA41;
  assign sine_lookup[208 ]    = 16'hFA7C;
  assign sine_lookup[209 ]    = 16'hFAB6;
  assign sine_lookup[210 ]    = 16'hFAEE;
  assign sine_lookup[211 ]    = 16'hFB26;
  assign sine_lookup[212 ]    = 16'hFB5C;
  assign sine_lookup[213 ]    = 16'hFB91;
  assign sine_lookup[214 ]    = 16'hFBC5;
  assign sine_lookup[215 ]    = 16'hFBF8;
  assign sine_lookup[216 ]    = 16'hFC29;
  assign sine_lookup[217 ]    = 16'hFC59;
  assign sine_lookup[218 ]    = 16'hFC88;
  assign sine_lookup[219 ]    = 16'hFCB6;
  assign sine_lookup[220 ]    = 16'hFCE3;
  assign sine_lookup[221 ]    = 16'hFD0E;
  assign sine_lookup[222 ]    = 16'hFD39;
  assign sine_lookup[223 ]    = 16'hFD62;
  assign sine_lookup[224 ]    = 16'hFD89;
  assign sine_lookup[225 ]    = 16'hFDB0;
  assign sine_lookup[226 ]    = 16'hFDD5;
  assign sine_lookup[227 ]    = 16'hFDFA;
  assign sine_lookup[228 ]    = 16'hFE1D;
  assign sine_lookup[229 ]    = 16'hFE3E;
  assign sine_lookup[230 ]    = 16'hFE5F;
  assign sine_lookup[231 ]    = 16'hFE7E;
  assign sine_lookup[232 ]    = 16'hFE9C;
  assign sine_lookup[233 ]    = 16'hFEB9;
  assign sine_lookup[234 ]    = 16'hFED5;
  assign sine_lookup[235 ]    = 16'hFEEF;
  assign sine_lookup[236 ]    = 16'hFF09;
  assign sine_lookup[237 ]    = 16'hFF21;
  assign sine_lookup[238 ]    = 16'hFF37;
  assign sine_lookup[239 ]    = 16'hFF4D;
  assign sine_lookup[240 ]    = 16'hFF61;
  assign sine_lookup[241 ]    = 16'hFF74;
  assign sine_lookup[242 ]    = 16'hFF86;
  assign sine_lookup[243 ]    = 16'hFF97;
  assign sine_lookup[244 ]    = 16'hFFA6;
  assign sine_lookup[245 ]    = 16'hFFB4;
  assign sine_lookup[246 ]    = 16'hFFC1;
  assign sine_lookup[247 ]    = 16'hFFCD;
  assign sine_lookup[248 ]    = 16'hFFD8;
  assign sine_lookup[249 ]    = 16'hFFE1;
  assign sine_lookup[250 ]    = 16'hFFE9;
  assign sine_lookup[251 ]    = 16'hFFF0;
  assign sine_lookup[252 ]    = 16'hFFF5;
  assign sine_lookup[253 ]    = 16'hFFF9;
  assign sine_lookup[254 ]    = 16'hFFFD;
  assign sine_lookup[255 ]    = 16'hFFFE;
  assign sine_lookup[256 ]    = 16'hFFFF;
  assign sine_lookup[257 ]    = 16'hFFFE;
  assign sine_lookup[258 ]    = 16'hFFFD;
  assign sine_lookup[259 ]    = 16'hFFF9;
  assign sine_lookup[260 ]    = 16'hFFF5;
  assign sine_lookup[261 ]    = 16'hFFF0;
  assign sine_lookup[262 ]    = 16'hFFE9;
  assign sine_lookup[263 ]    = 16'hFFE1;
  assign sine_lookup[264 ]    = 16'hFFD8;
  assign sine_lookup[265 ]    = 16'hFFCD;
  assign sine_lookup[266 ]    = 16'hFFC1;
  assign sine_lookup[267 ]    = 16'hFFB4;
  assign sine_lookup[268 ]    = 16'hFFA6;
  assign sine_lookup[269 ]    = 16'hFF97;
  assign sine_lookup[270 ]    = 16'hFF86;
  assign sine_lookup[271 ]    = 16'hFF74;
  assign sine_lookup[272 ]    = 16'hFF61;
  assign sine_lookup[273 ]    = 16'hFF4D;
  assign sine_lookup[274 ]    = 16'hFF37;
  assign sine_lookup[275 ]    = 16'hFF21;
  assign sine_lookup[276 ]    = 16'hFF09;
  assign sine_lookup[277 ]    = 16'hFEEF;
  assign sine_lookup[278 ]    = 16'hFED5;
  assign sine_lookup[279 ]    = 16'hFEB9;
  assign sine_lookup[280 ]    = 16'hFE9C;
  assign sine_lookup[281 ]    = 16'hFE7E;
  assign sine_lookup[282 ]    = 16'hFE5F;
  assign sine_lookup[283 ]    = 16'hFE3E;
  assign sine_lookup[284 ]    = 16'hFE1D;
  assign sine_lookup[285 ]    = 16'hFDFA;
  assign sine_lookup[286 ]    = 16'hFDD5;
  assign sine_lookup[287 ]    = 16'hFDB0;
  assign sine_lookup[288 ]    = 16'hFD89;
  assign sine_lookup[289 ]    = 16'hFD62;
  assign sine_lookup[290 ]    = 16'hFD39;
  assign sine_lookup[291 ]    = 16'hFD0E;
  assign sine_lookup[292 ]    = 16'hFCE3;
  assign sine_lookup[293 ]    = 16'hFCB6;
  assign sine_lookup[294 ]    = 16'hFC88;
  assign sine_lookup[295 ]    = 16'hFC59;
  assign sine_lookup[296 ]    = 16'hFC29;
  assign sine_lookup[297 ]    = 16'hFBF8;
  assign sine_lookup[298 ]    = 16'hFBC5;
  assign sine_lookup[299 ]    = 16'hFB91;
  assign sine_lookup[300 ]    = 16'hFB5C;
  assign sine_lookup[301 ]    = 16'hFB26;
  assign sine_lookup[302 ]    = 16'hFAEE;
  assign sine_lookup[303 ]    = 16'hFAB6;
  assign sine_lookup[304 ]    = 16'hFA7C;
  assign sine_lookup[305 ]    = 16'hFA41;
  assign sine_lookup[306 ]    = 16'hFA05;
  assign sine_lookup[307 ]    = 16'hF9C8;
  assign sine_lookup[308 ]    = 16'hF989;
  assign sine_lookup[309 ]    = 16'hF94A;
  assign sine_lookup[310 ]    = 16'hF909;
  assign sine_lookup[311 ]    = 16'hF8C7;
  assign sine_lookup[312 ]    = 16'hF884;
  assign sine_lookup[313 ]    = 16'hF83F;
  assign sine_lookup[314 ]    = 16'hF7FA;
  assign sine_lookup[315 ]    = 16'hF7B3;
  assign sine_lookup[316 ]    = 16'hF76B;
  assign sine_lookup[317 ]    = 16'hF722;
  assign sine_lookup[318 ]    = 16'hF6D8;
  assign sine_lookup[319 ]    = 16'hF68D;
  assign sine_lookup[320 ]    = 16'hF641;
  assign sine_lookup[321 ]    = 16'hF5F3;
  assign sine_lookup[322 ]    = 16'hF5A5;
  assign sine_lookup[323 ]    = 16'hF555;
  assign sine_lookup[324 ]    = 16'hF504;
  assign sine_lookup[325 ]    = 16'hF4B2;
  assign sine_lookup[326 ]    = 16'hF45F;
  assign sine_lookup[327 ]    = 16'hF40A;
  assign sine_lookup[328 ]    = 16'hF3B5;
  assign sine_lookup[329 ]    = 16'hF35E;
  assign sine_lookup[330 ]    = 16'hF307;
  assign sine_lookup[331 ]    = 16'hF2AE;
  assign sine_lookup[332 ]    = 16'hF254;
  assign sine_lookup[333 ]    = 16'hF1F9;
  assign sine_lookup[334 ]    = 16'hF19D;
  assign sine_lookup[335 ]    = 16'hF140;
  assign sine_lookup[336 ]    = 16'hF0E2;
  assign sine_lookup[337 ]    = 16'hF083;
  assign sine_lookup[338 ]    = 16'hF022;
  assign sine_lookup[339 ]    = 16'hEFC1;
  assign sine_lookup[340 ]    = 16'hEF5E;
  assign sine_lookup[341 ]    = 16'hEEFB;
  assign sine_lookup[342 ]    = 16'hEE96;
  assign sine_lookup[343 ]    = 16'hEE30;
  assign sine_lookup[344 ]    = 16'hEDC9;
  assign sine_lookup[345 ]    = 16'hED61;
  assign sine_lookup[346 ]    = 16'hECF8;
  assign sine_lookup[347 ]    = 16'hEC8E;
  assign sine_lookup[348 ]    = 16'hEC23;
  assign sine_lookup[349 ]    = 16'hEBB7;
  assign sine_lookup[350 ]    = 16'hEB4A;
  assign sine_lookup[351 ]    = 16'hEADC;
  assign sine_lookup[352 ]    = 16'hEA6D;
  assign sine_lookup[353 ]    = 16'hE9FD;
  assign sine_lookup[354 ]    = 16'hE98B;
  assign sine_lookup[355 ]    = 16'hE919;
  assign sine_lookup[356 ]    = 16'hE8A6;
  assign sine_lookup[357 ]    = 16'hE832;
  assign sine_lookup[358 ]    = 16'hE7BC;
  assign sine_lookup[359 ]    = 16'hE746;
  assign sine_lookup[360 ]    = 16'hE6CF;
  assign sine_lookup[361 ]    = 16'hE656;
  assign sine_lookup[362 ]    = 16'hE5DD;
  assign sine_lookup[363 ]    = 16'hE563;
  assign sine_lookup[364 ]    = 16'hE4E8;
  assign sine_lookup[365 ]    = 16'hE46C;
  assign sine_lookup[366 ]    = 16'hE3EE;
  assign sine_lookup[367 ]    = 16'hE370;
  assign sine_lookup[368 ]    = 16'hE2F1;
  assign sine_lookup[369 ]    = 16'hE271;
  assign sine_lookup[370 ]    = 16'hE1F0;
  assign sine_lookup[371 ]    = 16'hE16E;
  assign sine_lookup[372 ]    = 16'hE0EB;
  assign sine_lookup[373 ]    = 16'hE068;
  assign sine_lookup[374 ]    = 16'hDFE3;
  assign sine_lookup[375 ]    = 16'hDF5D;
  assign sine_lookup[376 ]    = 16'hDED7;
  assign sine_lookup[377 ]    = 16'hDE4F;
  assign sine_lookup[378 ]    = 16'hDDC7;
  assign sine_lookup[379 ]    = 16'hDD3E;
  assign sine_lookup[380 ]    = 16'hDCB3;
  assign sine_lookup[381 ]    = 16'hDC28;
  assign sine_lookup[382 ]    = 16'hDB9C;
  assign sine_lookup[383 ]    = 16'hDB0F;
  assign sine_lookup[384 ]    = 16'hDA82;
  assign sine_lookup[385 ]    = 16'hD9F3;
  assign sine_lookup[386 ]    = 16'hD964;
  assign sine_lookup[387 ]    = 16'hD8D3;
  assign sine_lookup[388 ]    = 16'hD842;
  assign sine_lookup[389 ]    = 16'hD7B0;
  assign sine_lookup[390 ]    = 16'hD71D;
  assign sine_lookup[391 ]    = 16'hD68A;
  assign sine_lookup[392 ]    = 16'hD5F5;
  assign sine_lookup[393 ]    = 16'hD560;
  assign sine_lookup[394 ]    = 16'hD4C9;
  assign sine_lookup[395 ]    = 16'hD432;
  assign sine_lookup[396 ]    = 16'hD39B;
  assign sine_lookup[397 ]    = 16'hD302;
  assign sine_lookup[398 ]    = 16'hD268;
  assign sine_lookup[399 ]    = 16'hD1CE;
  assign sine_lookup[400 ]    = 16'hD133;
  assign sine_lookup[401 ]    = 16'hD097;
  assign sine_lookup[402 ]    = 16'hCFFB;
  assign sine_lookup[403 ]    = 16'hCF5D;
  assign sine_lookup[404 ]    = 16'hCEBF;
  assign sine_lookup[405 ]    = 16'hCE20;
  assign sine_lookup[406 ]    = 16'hCD81;
  assign sine_lookup[407 ]    = 16'hCCE0;
  assign sine_lookup[408 ]    = 16'hCC3F;
  assign sine_lookup[409 ]    = 16'hCB9D;
  assign sine_lookup[410 ]    = 16'hCAFB;
  assign sine_lookup[411 ]    = 16'hCA58;
  assign sine_lookup[412 ]    = 16'hC9B4;
  assign sine_lookup[413 ]    = 16'hC90F;
  assign sine_lookup[414 ]    = 16'hC869;
  assign sine_lookup[415 ]    = 16'hC7C3;
  assign sine_lookup[416 ]    = 16'hC71C;
  assign sine_lookup[417 ]    = 16'hC675;
  assign sine_lookup[418 ]    = 16'hC5CD;
  assign sine_lookup[419 ]    = 16'hC524;
  assign sine_lookup[420 ]    = 16'hC47A;
  assign sine_lookup[421 ]    = 16'hC3D0;
  assign sine_lookup[422 ]    = 16'hC325;
  assign sine_lookup[423 ]    = 16'hC27A;
  assign sine_lookup[424 ]    = 16'hC1CE;
  assign sine_lookup[425 ]    = 16'hC121;
  assign sine_lookup[426 ]    = 16'hC073;
  assign sine_lookup[427 ]    = 16'hBFC5;
  assign sine_lookup[428 ]    = 16'hBF17;
  assign sine_lookup[429 ]    = 16'hBE68;
  assign sine_lookup[430 ]    = 16'hBDB8;
  assign sine_lookup[431 ]    = 16'hBD07;
  assign sine_lookup[432 ]    = 16'hBC56;
  assign sine_lookup[433 ]    = 16'hBBA5;
  assign sine_lookup[434 ]    = 16'hBAF2;
  assign sine_lookup[435 ]    = 16'hBA40;
  assign sine_lookup[436 ]    = 16'hB98C;
  assign sine_lookup[437 ]    = 16'hB8D9;
  assign sine_lookup[438 ]    = 16'hB824;
  assign sine_lookup[439 ]    = 16'hB76F;
  assign sine_lookup[440 ]    = 16'hB6BA;
  assign sine_lookup[441 ]    = 16'hB604;
  assign sine_lookup[442 ]    = 16'hB54D;
  assign sine_lookup[443 ]    = 16'hB496;
  assign sine_lookup[444 ]    = 16'hB3DF;
  assign sine_lookup[445 ]    = 16'hB326;
  assign sine_lookup[446 ]    = 16'hB26E;
  assign sine_lookup[447 ]    = 16'hB1B5;
  assign sine_lookup[448 ]    = 16'hB0FB;
  assign sine_lookup[449 ]    = 16'hB041;
  assign sine_lookup[450 ]    = 16'hAF87;
  assign sine_lookup[451 ]    = 16'hAECC;
  assign sine_lookup[452 ]    = 16'hAE11;
  assign sine_lookup[453 ]    = 16'hAD55;
  assign sine_lookup[454 ]    = 16'hAC99;
  assign sine_lookup[455 ]    = 16'hABDC;
  assign sine_lookup[456 ]    = 16'hAB1F;
  assign sine_lookup[457 ]    = 16'hAA61;
  assign sine_lookup[458 ]    = 16'hA9A3;
  assign sine_lookup[459 ]    = 16'hA8E5;
  assign sine_lookup[460 ]    = 16'hA826;
  assign sine_lookup[461 ]    = 16'hA767;
  assign sine_lookup[462 ]    = 16'hA6A8;
  assign sine_lookup[463 ]    = 16'hA5E8;
  assign sine_lookup[464 ]    = 16'hA528;
  assign sine_lookup[465 ]    = 16'hA467;
  assign sine_lookup[466 ]    = 16'hA3A6;
  assign sine_lookup[467 ]    = 16'hA2E5;
  assign sine_lookup[468 ]    = 16'hA223;
  assign sine_lookup[469 ]    = 16'hA161;
  assign sine_lookup[470 ]    = 16'hA09F;
  assign sine_lookup[471 ]    = 16'h9FDD;
  assign sine_lookup[472 ]    = 16'h9F1A;
  assign sine_lookup[473 ]    = 16'h9E57;
  assign sine_lookup[474 ]    = 16'h9D93;
  assign sine_lookup[475 ]    = 16'h9CCF;
  assign sine_lookup[476 ]    = 16'h9C0B;
  assign sine_lookup[477 ]    = 16'h9B47;
  assign sine_lookup[478 ]    = 16'h9A82;
  assign sine_lookup[479 ]    = 16'h99BE;
  assign sine_lookup[480 ]    = 16'h98F9;
  assign sine_lookup[481 ]    = 16'h9833;
  assign sine_lookup[482 ]    = 16'h976E;
  assign sine_lookup[483 ]    = 16'h96A8;
  assign sine_lookup[484 ]    = 16'h95E2;
  assign sine_lookup[485 ]    = 16'h951C;
  assign sine_lookup[486 ]    = 16'h9455;
  assign sine_lookup[487 ]    = 16'h938F;
  assign sine_lookup[488 ]    = 16'h92C8;
  assign sine_lookup[489 ]    = 16'h9201;
  assign sine_lookup[490 ]    = 16'h913A;
  assign sine_lookup[491 ]    = 16'h9072;
  assign sine_lookup[492 ]    = 16'h8FAB;
  assign sine_lookup[493 ]    = 16'h8EE3;
  assign sine_lookup[494 ]    = 16'h8E1C;
  assign sine_lookup[495 ]    = 16'h8D54;
  assign sine_lookup[496 ]    = 16'h8C8C;
  assign sine_lookup[497 ]    = 16'h8BC4;
  assign sine_lookup[498 ]    = 16'h8AFB;
  assign sine_lookup[499 ]    = 16'h8A33;
  assign sine_lookup[500 ]    = 16'h896A;
  assign sine_lookup[501 ]    = 16'h88A2;
  assign sine_lookup[502 ]    = 16'h87D9;
  assign sine_lookup[503 ]    = 16'h8711;
  assign sine_lookup[504 ]    = 16'h8648;
  assign sine_lookup[505 ]    = 16'h857F;
  assign sine_lookup[506 ]    = 16'h84B6;
  assign sine_lookup[507 ]    = 16'h83ED;
  assign sine_lookup[508 ]    = 16'h8324;
  assign sine_lookup[509 ]    = 16'h825B;
  assign sine_lookup[510 ]    = 16'h8192;
  assign sine_lookup[511 ]    = 16'h80C9;
  assign sine_lookup[512 ]    = 16'h8000;
  assign sine_lookup[513 ]    = 16'h7F37;
  assign sine_lookup[514 ]    = 16'h7E6E;
  assign sine_lookup[515 ]    = 16'h7DA5;
  assign sine_lookup[516 ]    = 16'h7CDC;
  assign sine_lookup[517 ]    = 16'h7C13;
  assign sine_lookup[518 ]    = 16'h7B4A;
  assign sine_lookup[519 ]    = 16'h7A81;
  assign sine_lookup[520 ]    = 16'h79B8;
  assign sine_lookup[521 ]    = 16'h78EF;
  assign sine_lookup[522 ]    = 16'h7827;
  assign sine_lookup[523 ]    = 16'h775E;
  assign sine_lookup[524 ]    = 16'h7696;
  assign sine_lookup[525 ]    = 16'h75CD;
  assign sine_lookup[526 ]    = 16'h7505;
  assign sine_lookup[527 ]    = 16'h743C;
  assign sine_lookup[528 ]    = 16'h7374;
  assign sine_lookup[529 ]    = 16'h72AC;
  assign sine_lookup[530 ]    = 16'h71E4;
  assign sine_lookup[531 ]    = 16'h711D;
  assign sine_lookup[532 ]    = 16'h7055;
  assign sine_lookup[533 ]    = 16'h6F8E;
  assign sine_lookup[534 ]    = 16'h6EC6;
  assign sine_lookup[535 ]    = 16'h6DFF;
  assign sine_lookup[536 ]    = 16'h6D38;
  assign sine_lookup[537 ]    = 16'h6C71;
  assign sine_lookup[538 ]    = 16'h6BAB;
  assign sine_lookup[539 ]    = 16'h6AE4;
  assign sine_lookup[540 ]    = 16'h6A1E;
  assign sine_lookup[541 ]    = 16'h6958;
  assign sine_lookup[542 ]    = 16'h6892;
  assign sine_lookup[543 ]    = 16'h67CD;
  assign sine_lookup[544 ]    = 16'h6707;
  assign sine_lookup[545 ]    = 16'h6642;
  assign sine_lookup[546 ]    = 16'h657E;
  assign sine_lookup[547 ]    = 16'h64B9;
  assign sine_lookup[548 ]    = 16'h63F5;
  assign sine_lookup[549 ]    = 16'h6331;
  assign sine_lookup[550 ]    = 16'h626D;
  assign sine_lookup[551 ]    = 16'h61A9;
  assign sine_lookup[552 ]    = 16'h60E6;
  assign sine_lookup[553 ]    = 16'h6023;
  assign sine_lookup[554 ]    = 16'h5F61;
  assign sine_lookup[555 ]    = 16'h5E9F;
  assign sine_lookup[556 ]    = 16'h5DDD;
  assign sine_lookup[557 ]    = 16'h5D1B;
  assign sine_lookup[558 ]    = 16'h5C5A;
  assign sine_lookup[559 ]    = 16'h5B99;
  assign sine_lookup[560 ]    = 16'h5AD8;
  assign sine_lookup[561 ]    = 16'h5A18;
  assign sine_lookup[562 ]    = 16'h5958;
  assign sine_lookup[563 ]    = 16'h5899;
  assign sine_lookup[564 ]    = 16'h57DA;
  assign sine_lookup[565 ]    = 16'h571B;
  assign sine_lookup[566 ]    = 16'h565D;
  assign sine_lookup[567 ]    = 16'h559F;
  assign sine_lookup[568 ]    = 16'h54E1;
  assign sine_lookup[569 ]    = 16'h5424;
  assign sine_lookup[570 ]    = 16'h5367;
  assign sine_lookup[571 ]    = 16'h52AB;
  assign sine_lookup[572 ]    = 16'h51EF;
  assign sine_lookup[573 ]    = 16'h5134;
  assign sine_lookup[574 ]    = 16'h5079;
  assign sine_lookup[575 ]    = 16'h4FBF;
  assign sine_lookup[576 ]    = 16'h4F05;
  assign sine_lookup[577 ]    = 16'h4E4B;
  assign sine_lookup[578 ]    = 16'h4D92;
  assign sine_lookup[579 ]    = 16'h4CDA;
  assign sine_lookup[580 ]    = 16'h4C21;
  assign sine_lookup[581 ]    = 16'h4B6A;
  assign sine_lookup[582 ]    = 16'h4AB3;
  assign sine_lookup[583 ]    = 16'h49FC;
  assign sine_lookup[584 ]    = 16'h4946;
  assign sine_lookup[585 ]    = 16'h4891;
  assign sine_lookup[586 ]    = 16'h47DC;
  assign sine_lookup[587 ]    = 16'h4727;
  assign sine_lookup[588 ]    = 16'h4674;
  assign sine_lookup[589 ]    = 16'h45C0;
  assign sine_lookup[590 ]    = 16'h450E;
  assign sine_lookup[591 ]    = 16'h445B;
  assign sine_lookup[592 ]    = 16'h43AA;
  assign sine_lookup[593 ]    = 16'h42F9;
  assign sine_lookup[594 ]    = 16'h4248;
  assign sine_lookup[595 ]    = 16'h4198;
  assign sine_lookup[596 ]    = 16'h40E9;
  assign sine_lookup[597 ]    = 16'h403B;
  assign sine_lookup[598 ]    = 16'h3F8D;
  assign sine_lookup[599 ]    = 16'h3EDF;
  assign sine_lookup[600 ]    = 16'h3E32;
  assign sine_lookup[601 ]    = 16'h3D86;
  assign sine_lookup[602 ]    = 16'h3CDB;
  assign sine_lookup[603 ]    = 16'h3C30;
  assign sine_lookup[604 ]    = 16'h3B86;
  assign sine_lookup[605 ]    = 16'h3ADC;
  assign sine_lookup[606 ]    = 16'h3A33;
  assign sine_lookup[607 ]    = 16'h398B;
  assign sine_lookup[608 ]    = 16'h38E4;
  assign sine_lookup[609 ]    = 16'h383D;
  assign sine_lookup[610 ]    = 16'h3797;
  assign sine_lookup[611 ]    = 16'h36F1;
  assign sine_lookup[612 ]    = 16'h364C;
  assign sine_lookup[613 ]    = 16'h35A8;
  assign sine_lookup[614 ]    = 16'h3505;
  assign sine_lookup[615 ]    = 16'h3463;
  assign sine_lookup[616 ]    = 16'h33C1;
  assign sine_lookup[617 ]    = 16'h3320;
  assign sine_lookup[618 ]    = 16'h327F;
  assign sine_lookup[619 ]    = 16'h31E0;
  assign sine_lookup[620 ]    = 16'h3141;
  assign sine_lookup[621 ]    = 16'h30A3;
  assign sine_lookup[622 ]    = 16'h3005;
  assign sine_lookup[623 ]    = 16'h2F69;
  assign sine_lookup[624 ]    = 16'h2ECD;
  assign sine_lookup[625 ]    = 16'h2E32;
  assign sine_lookup[626 ]    = 16'h2D98;
  assign sine_lookup[627 ]    = 16'h2CFE;
  assign sine_lookup[628 ]    = 16'h2C65;
  assign sine_lookup[629 ]    = 16'h2BCE;
  assign sine_lookup[630 ]    = 16'h2B37;
  assign sine_lookup[631 ]    = 16'h2AA0;
  assign sine_lookup[632 ]    = 16'h2A0B;
  assign sine_lookup[633 ]    = 16'h2976;
  assign sine_lookup[634 ]    = 16'h28E3;
  assign sine_lookup[635 ]    = 16'h2850;
  assign sine_lookup[636 ]    = 16'h27BE;
  assign sine_lookup[637 ]    = 16'h272D;
  assign sine_lookup[638 ]    = 16'h269C;
  assign sine_lookup[639 ]    = 16'h260D;
  assign sine_lookup[640 ]    = 16'h257E;
  assign sine_lookup[641 ]    = 16'h24F1;
  assign sine_lookup[642 ]    = 16'h2464;
  assign sine_lookup[643 ]    = 16'h23D8;
  assign sine_lookup[644 ]    = 16'h234D;
  assign sine_lookup[645 ]    = 16'h22C2;
  assign sine_lookup[646 ]    = 16'h2239;
  assign sine_lookup[647 ]    = 16'h21B1;
  assign sine_lookup[648 ]    = 16'h2129;
  assign sine_lookup[649 ]    = 16'h20A3;
  assign sine_lookup[650 ]    = 16'h201D;
  assign sine_lookup[651 ]    = 16'h1F98;
  assign sine_lookup[652 ]    = 16'h1F15;
  assign sine_lookup[653 ]    = 16'h1E92;
  assign sine_lookup[654 ]    = 16'h1E10;
  assign sine_lookup[655 ]    = 16'h1D8F;
  assign sine_lookup[656 ]    = 16'h1D0F;
  assign sine_lookup[657 ]    = 16'h1C90;
  assign sine_lookup[658 ]    = 16'h1C12;
  assign sine_lookup[659 ]    = 16'h1B94;
  assign sine_lookup[660 ]    = 16'h1B18;
  assign sine_lookup[661 ]    = 16'h1A9D;
  assign sine_lookup[662 ]    = 16'h1A23;
  assign sine_lookup[663 ]    = 16'h19AA;
  assign sine_lookup[664 ]    = 16'h1931;
  assign sine_lookup[665 ]    = 16'h18BA;
  assign sine_lookup[666 ]    = 16'h1844;
  assign sine_lookup[667 ]    = 16'h17CE;
  assign sine_lookup[668 ]    = 16'h175A;
  assign sine_lookup[669 ]    = 16'h16E7;
  assign sine_lookup[670 ]    = 16'h1675;
  assign sine_lookup[671 ]    = 16'h1603;
  assign sine_lookup[672 ]    = 16'h1593;
  assign sine_lookup[673 ]    = 16'h1524;
  assign sine_lookup[674 ]    = 16'h14B6;
  assign sine_lookup[675 ]    = 16'h1449;
  assign sine_lookup[676 ]    = 16'h13DD;
  assign sine_lookup[677 ]    = 16'h1372;
  assign sine_lookup[678 ]    = 16'h1308;
  assign sine_lookup[679 ]    = 16'h129F;
  assign sine_lookup[680 ]    = 16'h1237;
  assign sine_lookup[681 ]    = 16'h11D0;
  assign sine_lookup[682 ]    = 16'h116A;
  assign sine_lookup[683 ]    = 16'h1105;
  assign sine_lookup[684 ]    = 16'h10A2;
  assign sine_lookup[685 ]    = 16'h103F;
  assign sine_lookup[686 ]    = 16'hFDE ;
  assign sine_lookup[687 ]    = 16'hF7D ;
  assign sine_lookup[688 ]    = 16'hF1E ;
  assign sine_lookup[689 ]    = 16'hEC0 ;
  assign sine_lookup[690 ]    = 16'hE63 ;
  assign sine_lookup[691 ]    = 16'hE07 ;
  assign sine_lookup[692 ]    = 16'hDAC ;
  assign sine_lookup[693 ]    = 16'hD52 ;
  assign sine_lookup[694 ]    = 16'hCF9 ;
  assign sine_lookup[695 ]    = 16'hCA2 ;
  assign sine_lookup[696 ]    = 16'hC4B ;
  assign sine_lookup[697 ]    = 16'hBF6 ;
  assign sine_lookup[698 ]    = 16'hBA1 ;
  assign sine_lookup[699 ]    = 16'hB4E ;
  assign sine_lookup[700 ]    = 16'hAFC ;
  assign sine_lookup[701 ]    = 16'hAAB ;
  assign sine_lookup[702 ]    = 16'hA5B ;
  assign sine_lookup[703 ]    = 16'hA0D ;
  assign sine_lookup[704 ]    = 16'h9BF ;
  assign sine_lookup[705 ]    = 16'h973 ;
  assign sine_lookup[706 ]    = 16'h928 ;
  assign sine_lookup[707 ]    = 16'h8DE ;
  assign sine_lookup[708 ]    = 16'h895 ;
  assign sine_lookup[709 ]    = 16'h84D ;
  assign sine_lookup[710 ]    = 16'h806 ;
  assign sine_lookup[711 ]    = 16'h7C1 ;
  assign sine_lookup[712 ]    = 16'h77C ;
  assign sine_lookup[713 ]    = 16'h739 ;
  assign sine_lookup[714 ]    = 16'h6F7 ;
  assign sine_lookup[715 ]    = 16'h6B6 ;
  assign sine_lookup[716 ]    = 16'h677 ;
  assign sine_lookup[717 ]    = 16'h638 ;
  assign sine_lookup[718 ]    = 16'h5FB ;
  assign sine_lookup[719 ]    = 16'h5BF ;
  assign sine_lookup[720 ]    = 16'h584 ;
  assign sine_lookup[721 ]    = 16'h54A ;
  assign sine_lookup[722 ]    = 16'h512 ;
  assign sine_lookup[723 ]    = 16'h4DA ;
  assign sine_lookup[724 ]    = 16'h4A4 ;
  assign sine_lookup[725 ]    = 16'h46F ;
  assign sine_lookup[726 ]    = 16'h43B ;
  assign sine_lookup[727 ]    = 16'h408 ;
  assign sine_lookup[728 ]    = 16'h3D7 ;
  assign sine_lookup[729 ]    = 16'h3A7 ;
  assign sine_lookup[730 ]    = 16'h378 ;
  assign sine_lookup[731 ]    = 16'h34A ;
  assign sine_lookup[732 ]    = 16'h31D ;
  assign sine_lookup[733 ]    = 16'h2F2 ;
  assign sine_lookup[734 ]    = 16'h2C7 ;
  assign sine_lookup[735 ]    = 16'h29E ;
  assign sine_lookup[736 ]    = 16'h277 ;
  assign sine_lookup[737 ]    = 16'h250 ;
  assign sine_lookup[738 ]    = 16'h22B ;
  assign sine_lookup[739 ]    = 16'h206 ;
  assign sine_lookup[740 ]    = 16'h1E3 ;
  assign sine_lookup[741 ]    = 16'h1C2 ;
  assign sine_lookup[742 ]    = 16'h1A1 ;
  assign sine_lookup[743 ]    = 16'h182 ;
  assign sine_lookup[744 ]    = 16'h164 ;
  assign sine_lookup[745 ]    = 16'h147 ;
  assign sine_lookup[746 ]    = 16'h12B ;
  assign sine_lookup[747 ]    = 16'h111 ;
  assign sine_lookup[748 ]    = 16'hF7  ;
  assign sine_lookup[749 ]    = 16'hDF  ;
  assign sine_lookup[750 ]    = 16'hC9  ;
  assign sine_lookup[751 ]    = 16'hB3  ;
  assign sine_lookup[752 ]    = 16'h9F  ;
  assign sine_lookup[753 ]    = 16'h8C  ;
  assign sine_lookup[754 ]    = 16'h7A  ;
  assign sine_lookup[755 ]    = 16'h69  ;
  assign sine_lookup[756 ]    = 16'h5A  ;
  assign sine_lookup[757 ]    = 16'h4C  ;
  assign sine_lookup[758 ]    = 16'h3F  ;
  assign sine_lookup[759 ]    = 16'h33  ;
  assign sine_lookup[760 ]    = 16'h28  ;
  assign sine_lookup[761 ]    = 16'h1F  ;
  assign sine_lookup[762 ]    = 16'h17  ;
  assign sine_lookup[763 ]    = 16'h10  ;
  assign sine_lookup[764 ]    = 16'hB   ;
  assign sine_lookup[765 ]    = 16'h7   ;
  assign sine_lookup[766 ]    = 16'h3   ;
  assign sine_lookup[767 ]    = 16'h2   ;
  assign sine_lookup[768 ]    = 16'h1   ;
  assign sine_lookup[769 ]    = 16'h2   ;
  assign sine_lookup[770 ]    = 16'h3   ;
  assign sine_lookup[771 ]    = 16'h7   ;
  assign sine_lookup[772 ]    = 16'hB   ;
  assign sine_lookup[773 ]    = 16'h10  ;
  assign sine_lookup[774 ]    = 16'h17  ;
  assign sine_lookup[775 ]    = 16'h1F  ;
  assign sine_lookup[776 ]    = 16'h28  ;
  assign sine_lookup[777 ]    = 16'h33  ;
  assign sine_lookup[778 ]    = 16'h3F  ;
  assign sine_lookup[779 ]    = 16'h4C  ;
  assign sine_lookup[780 ]    = 16'h5A  ;
  assign sine_lookup[781 ]    = 16'h69  ;
  assign sine_lookup[782 ]    = 16'h7A  ;
  assign sine_lookup[783 ]    = 16'h8C  ;
  assign sine_lookup[784 ]    = 16'h9F  ;
  assign sine_lookup[785 ]    = 16'hB3  ;
  assign sine_lookup[786 ]    = 16'hC9  ;
  assign sine_lookup[787 ]    = 16'hDF  ;
  assign sine_lookup[788 ]    = 16'hF7  ;
  assign sine_lookup[789 ]    = 16'h111 ;
  assign sine_lookup[790 ]    = 16'h12B ;
  assign sine_lookup[791 ]    = 16'h147 ;
  assign sine_lookup[792 ]    = 16'h164 ;
  assign sine_lookup[793 ]    = 16'h182 ;
  assign sine_lookup[794 ]    = 16'h1A1 ;
  assign sine_lookup[795 ]    = 16'h1C2 ;
  assign sine_lookup[796 ]    = 16'h1E3 ;
  assign sine_lookup[797 ]    = 16'h206 ;
  assign sine_lookup[798 ]    = 16'h22B ;
  assign sine_lookup[799 ]    = 16'h250 ;
  assign sine_lookup[800 ]    = 16'h277 ;
  assign sine_lookup[801 ]    = 16'h29E ;
  assign sine_lookup[802 ]    = 16'h2C7 ;
  assign sine_lookup[803 ]    = 16'h2F2 ;
  assign sine_lookup[804 ]    = 16'h31D ;
  assign sine_lookup[805 ]    = 16'h34A ;
  assign sine_lookup[806 ]    = 16'h378 ;
  assign sine_lookup[807 ]    = 16'h3A7 ;
  assign sine_lookup[808 ]    = 16'h3D7 ;
  assign sine_lookup[809 ]    = 16'h408 ;
  assign sine_lookup[810 ]    = 16'h43B ;
  assign sine_lookup[811 ]    = 16'h46F ;
  assign sine_lookup[812 ]    = 16'h4A4 ;
  assign sine_lookup[813 ]    = 16'h4DA ;
  assign sine_lookup[814 ]    = 16'h512 ;
  assign sine_lookup[815 ]    = 16'h54A ;
  assign sine_lookup[816 ]    = 16'h584 ;
  assign sine_lookup[817 ]    = 16'h5BF ;
  assign sine_lookup[818 ]    = 16'h5FB ;
  assign sine_lookup[819 ]    = 16'h638 ;
  assign sine_lookup[820 ]    = 16'h677 ;
  assign sine_lookup[821 ]    = 16'h6B6 ;
  assign sine_lookup[822 ]    = 16'h6F7 ;
  assign sine_lookup[823 ]    = 16'h739 ;
  assign sine_lookup[824 ]    = 16'h77C ;
  assign sine_lookup[825 ]    = 16'h7C1 ;
  assign sine_lookup[826 ]    = 16'h806 ;
  assign sine_lookup[827 ]    = 16'h84D ;
  assign sine_lookup[828 ]    = 16'h895 ;
  assign sine_lookup[829 ]    = 16'h8DE ;
  assign sine_lookup[830 ]    = 16'h928 ;
  assign sine_lookup[831 ]    = 16'h973 ;
  assign sine_lookup[832 ]    = 16'h9BF ;
  assign sine_lookup[833 ]    = 16'hA0D ;
  assign sine_lookup[834 ]    = 16'hA5B ;
  assign sine_lookup[835 ]    = 16'hAAB ;
  assign sine_lookup[836 ]    = 16'hAFC ;
  assign sine_lookup[837 ]    = 16'hB4E ;
  assign sine_lookup[838 ]    = 16'hBA1 ;
  assign sine_lookup[839 ]    = 16'hBF6 ;
  assign sine_lookup[840 ]    = 16'hC4B ;
  assign sine_lookup[841 ]    = 16'hCA2 ;
  assign sine_lookup[842 ]    = 16'hCF9 ;
  assign sine_lookup[843 ]    = 16'hD52 ;
  assign sine_lookup[844 ]    = 16'hDAC ;
  assign sine_lookup[845 ]    = 16'hE07 ;
  assign sine_lookup[846 ]    = 16'hE63 ;
  assign sine_lookup[847 ]    = 16'hEC0 ;
  assign sine_lookup[848 ]    = 16'hF1E ;
  assign sine_lookup[849 ]    = 16'hF7D ;
  assign sine_lookup[850 ]    = 16'hFDE ;
  assign sine_lookup[851 ]    = 16'h103F;
  assign sine_lookup[852 ]    = 16'h10A2;
  assign sine_lookup[853 ]    = 16'h1105;
  assign sine_lookup[854 ]    = 16'h116A;
  assign sine_lookup[855 ]    = 16'h11D0;
  assign sine_lookup[856 ]    = 16'h1237;
  assign sine_lookup[857 ]    = 16'h129F;
  assign sine_lookup[858 ]    = 16'h1308;
  assign sine_lookup[859 ]    = 16'h1372;
  assign sine_lookup[860 ]    = 16'h13DD;
  assign sine_lookup[861 ]    = 16'h1449;
  assign sine_lookup[862 ]    = 16'h14B6;
  assign sine_lookup[863 ]    = 16'h1524;
  assign sine_lookup[864 ]    = 16'h1593;
  assign sine_lookup[865 ]    = 16'h1603;
  assign sine_lookup[866 ]    = 16'h1675;
  assign sine_lookup[867 ]    = 16'h16E7;
  assign sine_lookup[868 ]    = 16'h175A;
  assign sine_lookup[869 ]    = 16'h17CE;
  assign sine_lookup[870 ]    = 16'h1844;
  assign sine_lookup[871 ]    = 16'h18BA;
  assign sine_lookup[872 ]    = 16'h1931;
  assign sine_lookup[873 ]    = 16'h19AA;
  assign sine_lookup[874 ]    = 16'h1A23;
  assign sine_lookup[875 ]    = 16'h1A9D;
  assign sine_lookup[876 ]    = 16'h1B18;
  assign sine_lookup[877 ]    = 16'h1B94;
  assign sine_lookup[878 ]    = 16'h1C12;
  assign sine_lookup[879 ]    = 16'h1C90;
  assign sine_lookup[880 ]    = 16'h1D0F;
  assign sine_lookup[881 ]    = 16'h1D8F;
  assign sine_lookup[882 ]    = 16'h1E10;
  assign sine_lookup[883 ]    = 16'h1E92;
  assign sine_lookup[884 ]    = 16'h1F15;
  assign sine_lookup[885 ]    = 16'h1F98;
  assign sine_lookup[886 ]    = 16'h201D;
  assign sine_lookup[887 ]    = 16'h20A3;
  assign sine_lookup[888 ]    = 16'h2129;
  assign sine_lookup[889 ]    = 16'h21B1;
  assign sine_lookup[890 ]    = 16'h2239;
  assign sine_lookup[891 ]    = 16'h22C2;
  assign sine_lookup[892 ]    = 16'h234D;
  assign sine_lookup[893 ]    = 16'h23D8;
  assign sine_lookup[894 ]    = 16'h2464;
  assign sine_lookup[895 ]    = 16'h24F1;
  assign sine_lookup[896 ]    = 16'h257E;
  assign sine_lookup[897 ]    = 16'h260D;
  assign sine_lookup[898 ]    = 16'h269C;
  assign sine_lookup[899 ]    = 16'h272D;
  assign sine_lookup[900 ]    = 16'h27BE;
  assign sine_lookup[901 ]    = 16'h2850;
  assign sine_lookup[902 ]    = 16'h28E3;
  assign sine_lookup[903 ]    = 16'h2976;
  assign sine_lookup[904 ]    = 16'h2A0B;
  assign sine_lookup[905 ]    = 16'h2AA0;
  assign sine_lookup[906 ]    = 16'h2B37;
  assign sine_lookup[907 ]    = 16'h2BCE;
  assign sine_lookup[908 ]    = 16'h2C65;
  assign sine_lookup[909 ]    = 16'h2CFE;
  assign sine_lookup[910 ]    = 16'h2D98;
  assign sine_lookup[911 ]    = 16'h2E32;
  assign sine_lookup[912 ]    = 16'h2ECD;
  assign sine_lookup[913 ]    = 16'h2F69;
  assign sine_lookup[914 ]    = 16'h3005;
  assign sine_lookup[915 ]    = 16'h30A3;
  assign sine_lookup[916 ]    = 16'h3141;
  assign sine_lookup[917 ]    = 16'h31E0;
  assign sine_lookup[918 ]    = 16'h327F;
  assign sine_lookup[919 ]    = 16'h3320;
  assign sine_lookup[920 ]    = 16'h33C1;
  assign sine_lookup[921 ]    = 16'h3463;
  assign sine_lookup[922 ]    = 16'h3505;
  assign sine_lookup[923 ]    = 16'h35A8;
  assign sine_lookup[924 ]    = 16'h364C;
  assign sine_lookup[925 ]    = 16'h36F1;
  assign sine_lookup[926 ]    = 16'h3797;
  assign sine_lookup[927 ]    = 16'h383D;
  assign sine_lookup[928 ]    = 16'h38E4;
  assign sine_lookup[929 ]    = 16'h398B;
  assign sine_lookup[930 ]    = 16'h3A33;
  assign sine_lookup[931 ]    = 16'h3ADC;
  assign sine_lookup[932 ]    = 16'h3B86;
  assign sine_lookup[933 ]    = 16'h3C30;
  assign sine_lookup[934 ]    = 16'h3CDB;
  assign sine_lookup[935 ]    = 16'h3D86;
  assign sine_lookup[936 ]    = 16'h3E32;
  assign sine_lookup[937 ]    = 16'h3EDF;
  assign sine_lookup[938 ]    = 16'h3F8D;
  assign sine_lookup[939 ]    = 16'h403B;
  assign sine_lookup[940 ]    = 16'h40E9;
  assign sine_lookup[941 ]    = 16'h4198;
  assign sine_lookup[942 ]    = 16'h4248;
  assign sine_lookup[943 ]    = 16'h42F9;
  assign sine_lookup[944 ]    = 16'h43AA;
  assign sine_lookup[945 ]    = 16'h445B;
  assign sine_lookup[946 ]    = 16'h450E;
  assign sine_lookup[947 ]    = 16'h45C0;
  assign sine_lookup[948 ]    = 16'h4674;
  assign sine_lookup[949 ]    = 16'h4727;
  assign sine_lookup[950 ]    = 16'h47DC;
  assign sine_lookup[951 ]    = 16'h4891;
  assign sine_lookup[952 ]    = 16'h4946;
  assign sine_lookup[953 ]    = 16'h49FC;
  assign sine_lookup[954 ]    = 16'h4AB3;
  assign sine_lookup[955 ]    = 16'h4B6A;
  assign sine_lookup[956 ]    = 16'h4C21;
  assign sine_lookup[957 ]    = 16'h4CDA;
  assign sine_lookup[958 ]    = 16'h4D92;
  assign sine_lookup[959 ]    = 16'h4E4B;
  assign sine_lookup[960 ]    = 16'h4F05;
  assign sine_lookup[961 ]    = 16'h4FBF;
  assign sine_lookup[962 ]    = 16'h5079;
  assign sine_lookup[963 ]    = 16'h5134;
  assign sine_lookup[964 ]    = 16'h51EF;
  assign sine_lookup[965 ]    = 16'h52AB;
  assign sine_lookup[966 ]    = 16'h5367;
  assign sine_lookup[967 ]    = 16'h5424;
  assign sine_lookup[968 ]    = 16'h54E1;
  assign sine_lookup[969 ]    = 16'h559F;
  assign sine_lookup[970 ]    = 16'h565D;
  assign sine_lookup[971 ]    = 16'h571B;
  assign sine_lookup[972 ]    = 16'h57DA;
  assign sine_lookup[973 ]    = 16'h5899;
  assign sine_lookup[974 ]    = 16'h5958;
  assign sine_lookup[975 ]    = 16'h5A18;
  assign sine_lookup[976 ]    = 16'h5AD8;
  assign sine_lookup[977 ]    = 16'h5B99;
  assign sine_lookup[978 ]    = 16'h5C5A;
  assign sine_lookup[979 ]    = 16'h5D1B;
  assign sine_lookup[980 ]    = 16'h5DDD;
  assign sine_lookup[981 ]    = 16'h5E9F;
  assign sine_lookup[982 ]    = 16'h5F61;
  assign sine_lookup[983 ]    = 16'h6023;
  assign sine_lookup[984 ]    = 16'h60E6;
  assign sine_lookup[985 ]    = 16'h61A9;
  assign sine_lookup[986 ]    = 16'h626D;
  assign sine_lookup[987 ]    = 16'h6331;
  assign sine_lookup[988 ]    = 16'h63F5;
  assign sine_lookup[989 ]    = 16'h64B9;
  assign sine_lookup[990 ]    = 16'h657E;
  assign sine_lookup[991 ]    = 16'h6642;
  assign sine_lookup[992 ]    = 16'h6707;
  assign sine_lookup[993 ]    = 16'h67CD;
  assign sine_lookup[994 ]    = 16'h6892;
  assign sine_lookup[995 ]    = 16'h6958;
  assign sine_lookup[996 ]    = 16'h6A1E;
  assign sine_lookup[997 ]    = 16'h6AE4;
  assign sine_lookup[998 ]    = 16'h6BAB;
  assign sine_lookup[999 ]    = 16'h6C71;
  assign sine_lookup[1000]    = 16'h6D38;
  assign sine_lookup[1001]    = 16'h6DFF;
  assign sine_lookup[1002]    = 16'h6EC6;
  assign sine_lookup[1003]    = 16'h6F8E;
  assign sine_lookup[1004]    = 16'h7055;
  assign sine_lookup[1005]    = 16'h711D;
  assign sine_lookup[1006]    = 16'h71E4;
  assign sine_lookup[1007]    = 16'h72AC;
  assign sine_lookup[1008]    = 16'h7374;
  assign sine_lookup[1009]    = 16'h743C;
  assign sine_lookup[1010]    = 16'h7505;
  assign sine_lookup[1011]    = 16'h75CD;
  assign sine_lookup[1012]    = 16'h7696;
  assign sine_lookup[1013]    = 16'h775E;
  assign sine_lookup[1014]    = 16'h7827;
  assign sine_lookup[1015]    = 16'h78EF;
  assign sine_lookup[1016]    = 16'h79B8;
  assign sine_lookup[1017]    = 16'h7A81;
  assign sine_lookup[1018]    = 16'h7B4A;
  assign sine_lookup[1019]    = 16'h7C13;
  assign sine_lookup[1020]    = 16'h7CDC;
  assign sine_lookup[1021]    = 16'h7DA5;
  assign sine_lookup[1022]    = 16'h7E6E;
  assign sine_lookup[1023]    = 16'h7F37;
